module vraklib

struct VRakLib {

}
