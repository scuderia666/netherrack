module net

pub struct Network {
}

pub fn (mut n Network) start() {
    println("hi")
}