module netherrack

pub struct Netherrack {
}

pub fn (mut n Netherrack) start() {
}
